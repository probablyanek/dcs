* 0;Circuit1.sph
**************************************************************************************************
*                                            Circuit Design netlist                                      *
*                             created by Ansys Electronics Desktop                            *
**************************************************************************************************

.option PARHIER='local'
.option max_messages=1

* begin toplevel circuit


.SUB Substrate MS( H=0.0016 Er=4.4 TAND=0 TANM=0 MSat=0 MRem=0 HU=0.025
+MET1=1.724138 T1=1.778e-05)

A1 Port1 Port2 W=0.00159089 P=0.0139828 COMPONENT=TRL SUBSTRATE=Substrate
A4 Port2 net_3 W=0.00159089 P=0.0139828 COMPONENT=TRL SUBSTRATE=Substrate
A8 Port3 Port4 W=0.00159089 P=0.0139828 COMPONENT=TRL SUBSTRATE=Substrate
A9 Port4 net_6 W=0.00159089 P=0.0139828 COMPONENT=TRL SUBSTRATE=Substrate
A12 net_6 net_3 W=0.00159089 P=0.0139828 COMPONENT=TRL SUBSTRATE=Substrate
A15 Port3 Port1 W=0.00159089 P=0.0139828 COMPONENT=TRL SUBSTRATE=Substrate
RPort1 Port1 0 PORTNUM=1 RZ=50 IZ=0 
.PORT Port1 0 1 RPort1 
RPort2 Port2 0 PORTNUM=2 RZ=50 IZ=0 
.PORT Port2 0 2 RPort2 
RPort3 Port3 0 PORTNUM=3 RZ=50 IZ=0 
.PORT Port3 0 3 RPort3 
RPort4 Port4 0 PORTNUM=4 RZ=50 IZ=0 
.PORT Port4 0 4 RPort4 

* end toplevel circuit
.LNA
+ LIN 401 1000000000 5000000000
+ FLAG='LNA'

.end
